`timescale 1ns/1ns

module AND(
    input a,   
    input b,    
    output out  
);
    assign out = a & b; 
endmodule

